`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    14:32:01 05/19/2018 
// Design Name: 
// Module Name:    buf8 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module buf8( 
       input [7:0] din, 
       output [7:0] dout 
    ); 
      assign dout = din; 
    endmodule

